----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:47:44 12/14/2014 
-- Design Name: 
-- Module Name:    ball_sprite - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.ALL;

entity ball_sprite is
	port
	(
		x : in STD_LOGIC_VECTOR(9 downto 0);
		colour	:	out STD_LOGIC_VECTOR(1 downto 0)
	);
end ball_sprite;

architecture Behavioral of ball_sprite is
type SPRITE_ROM is array(integer range <>) of STD_LOGIC_VECTOR(1 downto 0);
constant rom : SPRITE_ROM (0 to 1023) := 
(	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,GREY_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	BLACK_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,GREY_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	BLACK_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,GREY_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	BLACK_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	GREY_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	GREY_2,GREY_2,GREY_2,BLACK_2,GREY_2,GREY_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,GREY_2,GREY_2,BLACK_2,GREY_2,GREY_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,BLACK_2,BLACK_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,GREY_2,GREY_2,GREY_2,GREY_2,WHITE_2,WHITE_2,WHITE_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,
	ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2,ALPHA_2);
begin
	colour <= rom(to_integer(unsigned(x)));
end Behavioral;

