----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:56:01 12/07/2014 
-- Design Name: 
-- Module Name:    cards_sprite - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cards_sprite_2 is
port
	(
		sprite_num	:	in		UNSIGNED(2 downto 0);
		x				:	in		STD_LOGIC_VECTOR(9 downto 0);
		draw_sprite	:	out	STD_LOGIC;
		rgb			:	out	STD_LOGIC_VECTOR(8 downto 0)
	);
end cards_sprite_2;

architecture Behavioral of cards_sprite_2 is
type CARDS_PALETTE is (BLACK, LIGHT_BLUE, WHITE, ORANGE, DARK_YELLOW, YELLOW, ALPHA);
type SPRITE_ROM is array (integer range <>) of CARDS_PALETTE;
constant BLACK_9 : std_logic_vector(8 downto 0) := "000000000";
constant LIGHT_BLUE_9 : std_logic_vector(8 downto 0) := "000100110";
constant WHITE_9 : std_logic_vector(8 downto 0) := "111111111";
constant ORANGE_9 : std_logic_vector(8 downto 0) := "111011001";
constant DARK_YELLOW_9 : std_logic_vector(8 downto 0) := "111101000";
constant YELLOW_9 : std_logic_vector(8 downto 0) := "111110000";
constant c_width : integer := 32;
constant c_height : integer := 32;
constant sprite_c4 : SPRITE_ROM (0 to 1023) := 
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,BLACK,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,ORANGE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,YELLOW,WHITE,BLACK,
BLACK,WHITE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,
BLACK,BLACK,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

constant sprite_c3 : SPRITE_ROM (0 to 1023) :=
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,DARK_YELLOW,DARK_YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,ORANGE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,ORANGE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,ORANGE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,YELLOW,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,YELLOW,LIGHT_BLUE,YELLOW,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,DARK_YELLOW,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,YELLOW,YELLOW,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,LIGHT_BLUE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

constant sprite_c2 : SPRITE_ROM (0 to 1023) :=
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,WHITE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);
constant sprite_c1 : SPRITE_ROM (0 to 1023) :=
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

signal rgb_dec,rgb_dec_4, rgb_dec_3, rgb_dec_2, rgb_dec_1  : CARDS_PALETTE;
begin
rgb_dec_4 <=	sprite_c4(to_integer(unsigned(x)));
rgb_dec_3 <=	sprite_c3(to_integer(unsigned(x)));
rgb_dec_2 <=	sprite_c2(to_integer(unsigned(x)));
rgb_dec_1 <=	sprite_c1(to_integer(unsigned(x)));
rgb_dec <=	rgb_dec_4 when sprite_num = 4 else
				rgb_dec_3 when sprite_num = 3 else
				rgb_dec_2 when sprite_num = 2 else
				rgb_dec_1 when sprite_num = 1 else
				ALPHA;
draw_sprite <= '1' when sprite_num /= 0 and rgb_dec /= ALPHA else '0';
rgb <=	WHITE_9 when rgb_dec = WHITE else
			LIGHT_BLUE_9 when rgb_dec = LIGHT_BLUE else
			ORANGE_9 when rgb_dec = ORANGE else
			DARK_YELLOW_9 when rgb_dec = DARK_YELLOW else
			YELLOW_9 when rgb_dec = YELLOW else
			BLACK_9;

end Behavioral;
