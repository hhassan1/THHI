----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:02:39 12/13/2014 
-- Design Name: 
-- Module Name:    moving_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.Types.ALL;

entity player_sprite_moving_1 is
	port
	(
		x : in STD_LOGIC_VECTOR(9 downto 0);
		colour	:	out STD_LOGIC_VECTOR(2 downto 0)
	);
end player_sprite_moving_1;

architecture Behavioral of player_sprite_moving_1 is
type SPRITE_ROM is array(integer range <>) of STD_LOGIC_VECTOR(2 downto 0);
constant rom : SPRITE_ROM(0 to 1023) :=
	(	ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,DARK_GREY_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,BLACK_3,DARK_RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,BLACK_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,WHITE_3,BLACK_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,
		BLACK_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,WHITE_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,BLACK_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,DARK_RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,
		BLACK_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,BLACK_3,ALPHA_3,ALPHA_3,
		BLACK_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,WHITE_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,RED_3,RED_3,RED_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,
		BLACK_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,
		BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,ALPHA_3,ALPHA_3,
		ALPHA_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,BLACK_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,WHITE_3,BLACK_3,ALPHA_3,ALPHA_3,
		ALPHA_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,DARK_GREY_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,SKIN_3,SKIN_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,BLACK_3,SKIN_3,SKIN_3,SKIN_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,WHITE_3,SKIN_3,BLACK_3,BLACK_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,BLACK_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,SKIN_3,SKIN_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,WHITE_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,BLACK_3,DARK_GREY_3,WHITE_3,WHITE_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,WHITE_3,WHITE_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,DARK_GREY_3,WHITE_3,WHITE_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,DARK_GREY_3,DARK_GREY_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,RED_3,RED_3,RED_3,RED_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,
		ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,BLACK_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3,ALPHA_3);
begin
	colour <= rom(to_integer(unsigned(x)));
end Behavioral;

