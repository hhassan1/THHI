----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:15:49 03/13/2015 
-- Design Name: 
-- Module Name:    endscreen - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity endscreen is
	port
	(
		win		:	in STD_LOGIC;
		vga_x		:	in UNSIGNED(9 downto 0);
		vga_y		:	in UNSIGNED(9 downto 0);
		draw_sprite	:	out STD_LOGIC
	);
end endscreen;

architecture Behavioral of endscreen is
type END_ROM is array(0 to 203) of STD_LOGIC;
constant win_rom : END_ROM := (
'1','0','0','0','1','0','0','1','1','0','0','1','0','0','1','0','1','0','0','1','0','0','1','0','1','0','1','0','0','0','1','0','0','0',
'0','1','0','1','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','1','0','0','1','0','0','0','1','1','0','0','1','0','0','0',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','1','0','0','1','0','1','0','1','0','1','0','1','0','0','0',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','1','0','0','1','0','1','0','1','0','0','1','1','0','0','0',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','1','0','0','1','0','1','0','1','0','0','0','1','0','0','0',
'0','0','1','0','0','0','0','1','1','0','0','0','1','1','0','0','0','1','1','0','1','1','0','0','1','0','1','0','0','0','1','0','0','0');
constant lose_rom : END_ROM := (
'1','0','0','0','1','0','0','1','1','0','0','1','0','0','1','0','1','0','0','0','0','1','1','0','0','0','1','1','1','0','1','1','1','1',
'0','1','0','1','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','0','1','0','0','1','0','1','0','0','0','0','1','0','0','0',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','0','1','0','0','1','0','1','1','1','0','0','1','1','1','1',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','0','1','0','0','1','0','0','0','0','1','0','1','0','0','0',
'0','0','1','0','0','0','1','0','0','1','0','1','0','0','1','0','1','0','0','0','1','0','0','1','0','0','0','0','1','0','1','0','0','0',
'0','0','1','0','0','0','0','1','1','0','0','0','1','1','0','0','1','1','1','0','0','1','1','0','0','1','1','1','0','0','1','1','1','1');
signal draw_win, draw_lose : STD_LOGIC;
begin
draw_win <= win_rom(to_integer(vga_x(9 downto 3) - 23 + (unsigned(std_logic_vector(vga_y(9 downto 3) - 27) & "00000")) + (unsigned(std_logic_vector(vga_y(9 downto 3) - 27) & "0"))));
draw_lose <= lose_rom(to_integer(vga_x(9 downto 3) - 23 + (unsigned(std_logic_vector(vga_y(9 downto 3) - 27) & "00000")) + (unsigned(std_logic_vector(vga_y(9 downto 3) - 27) & "0"))));
draw_sprite <= '0' when vga_x(9 downto 3) < 23 or vga_x(9 downto 3) >= 57 or vga_y(9 downto 3) < 27 or vga_y(9 downto 3) >= 33 else
					draw_win when win = '1' else
					draw_lose;
end Behavioral;

