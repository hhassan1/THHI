----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:56:01 12/07/2014 
-- Design Name: 
-- Module Name:    cards_sprite - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cards_sprite_3 is
port
	(
		sprite_num	:	in		UNSIGNED(2 downto 0);
		x				:	in		STD_LOGIC_VECTOR(9 downto 0);
		draw_sprite	:	out	STD_LOGIC;
		rgb			:	out	STD_LOGIC_VECTOR(8 downto 0)
	);
end cards_sprite_3;

architecture Behavioral of cards_sprite_3 is
type CARDS_PALETTE is (BLACK, BLUE_GREY, LIGHT_GREEN, LIME, PURPLE, DARK_GREEN, GREEN, BLUE, ALPHA);
type SPRITE_ROM is array (integer range <>) of CARDS_PALETTE;
constant BLACK_9 : std_logic_vector(8 downto 0) := "000000000";
constant BLUE_GREY_9 : std_logic_vector(8 downto 0) := "011100101";
constant LIGHT_GREEN_9 : std_logic_vector(8 downto 0) := "000111011";
constant LIME_9 : std_logic_vector(8 downto 0) := "011111011";
constant PURPLE_9 : std_logic_vector(8 downto 0) := "001001101";
constant DARK_GREEN_9 : std_logic_vector(8 downto 0) := "000011001";
constant GREEN_9 : std_logic_vector(8 downto 0) := "000100010";
constant BLUE_9 : std_logic_vector(8 downto 0) := "000000111";
constant c_width : integer := 32;
constant c_height : integer := 32;
constant sprite_c4 : SPRITE_ROM (0 to 1023) := 
(BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,PURPLE,PURPLE,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,PURPLE,PURPLE,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,LIME,LIGHT_GREEN,PURPLE,PURPLE,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,PURPLE,PURPLE,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,LIME,LIGHT_GREEN,LIME,PURPLE,PURPLE,LIGHT_GREEN,LIME,BLUE_GREY,BLUE_GREY,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,BLACK,
BLACK,LIGHT_GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,LIGHT_GREEN,BLUE,BLUE,BLUE,BLUE,GREEN,LIGHT_GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,BLUE,BLUE,BLUE,BLUE,GREEN,GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,LIGHT_GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,LIGHT_GREEN,BLUE,BLUE,LIGHT_GREEN,GREEN,GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,LIGHT_GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,LIGHT_GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLUE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,BLUE,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,BLUE,BLUE,GREEN,GREEN,BLUE,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,BLUE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,GREEN,BLUE,GREEN,GREEN,GREEN,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,BLUE,BLUE,BLUE,BLUE,BLUE,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,BLUE,BLUE,BLUE,BLUE,BLUE,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,BLUE,BLUE,BLUE,GREEN,GREEN,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,BLUE,BLUE,BLUE,GREEN,GREEN,BLUE,BLUE,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLACK,GREEN,GREEN,GREEN,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,GREEN,GREEN,GREEN,BLACK,
BLUE_GREY,BLUE_GREY,DARK_GREEN,DARK_GREEN,PURPLE,PURPLE,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,PURPLE,PURPLE,GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,DARK_GREEN,GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,
BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLUE_GREY);

constant sprite_c3 : SPRITE_ROM (0 to 1023) := 
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,LIME,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,LIME,LIME,LIME,LIME,LIME,LIME,PURPLE,LIME,LIME,LIME,LIME,LIME,LIME,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,LIGHT_GREEN,LIME,LIGHT_GREEN,LIME,LIGHT_GREEN,LIME,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIME,LIGHT_GREEN,LIME,LIGHT_GREEN,LIME,LIGHT_GREEN,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,LIGHT_GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,PURPLE,PURPLE,PURPLE,LIGHT_GREEN,PURPLE,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,LIGHT_GREEN,GREEN,PURPLE,GREEN,LIGHT_GREEN,PURPLE,LIGHT_GREEN,GREEN,PURPLE,LIGHT_GREEN,GREEN,PURPLE,PURPLE,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,PURPLE,PURPLE,GREEN,GREEN,PURPLE,GREEN,PURPLE,PURPLE,PURPLE,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,PURPLE,GREEN,PURPLE,GREEN,PURPLE,GREEN,PURPLE,PURPLE,PURPLE,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,PURPLE,PURPLE,PURPLE,GREEN,PURPLE,GREEN,PURPLE,PURPLE,PURPLE,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,GREEN,GREEN,GREEN,GREEN,GREEN,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,PURPLE,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,DARK_GREEN,PURPLE,DARK_GREEN,GREEN,DARK_GREEN,GREEN,DARK_GREEN,GREEN,DARK_GREEN,GREEN,DARK_GREEN,GREEN,DARK_GREEN,PURPLE,DARK_GREEN,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,DARK_GREEN,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLUE_GREY,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

constant sprite_c2 : SPRITE_ROM (0 to 1023) :=
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,LIGHT_GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,GREEN,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLUE_GREY,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

constant sprite_c1 : SPRITE_ROM (0 to 1023) :=
(BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,ALPHA,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,
BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK,BLACK);

signal rgb_dec,rgb_dec_4, rgb_dec_3, rgb_dec_2, rgb_dec_1  : CARDS_PALETTE;
begin
rgb_dec_4 <=	sprite_c4(to_integer(unsigned(x)));
rgb_dec_3 <=	sprite_c3(to_integer(unsigned(x)));
rgb_dec_2 <=	sprite_c2(to_integer(unsigned(x)));
rgb_dec_1 <=	sprite_c1(to_integer(unsigned(x)));
rgb_dec <=	rgb_dec_4 when sprite_num = 4 else
				rgb_dec_3 when sprite_num = 3 else
				rgb_dec_2 when sprite_num = 2 else
				rgb_dec_1 when sprite_num = 1 else
				ALPHA;
draw_sprite <= '1' when sprite_num /= 0 and rgb_dec /= ALPHA else '0';

rgb <=	BLUE_GREY_9 when rgb_dec = BLUE_GREY else
			BLUE_9 when rgb_dec = BLUE else
			LIGHT_GREEN_9 when rgb_dec = LIGHT_GREEN else
			GREEN_9 when rgb_dec = GREEN else
			DARK_GREEN_9 when rgb_dec = DARK_GREEN else
			PURPLE_9 when rgb_dec = PURPLE else
			LIME_9 when rgb_dec = LIME else
			BLACK_9;


end Behavioral;
